module clock_tree ( clk, 
  sink0,
  sink1,
  sink2,
  sink3,
  sink4,
  sink5,
  sink6,
  sink7,
  sink8,
  sink9,
  sink10,
  sink11,
  sink12,
  sink13,
  sink14,
  sink15,
  sink16,
  sink17,
  sink18,
  sink19,
  sink20,
  sink21,
  sink22,
  sink23,
  sink24,
  sink25,
  sink26,
  sink27,
  sink28,
  sink29,
  sink30,
  sink31,
  sink32,
  sink33,
  sink34,
  sink35,
  sink36,
  sink37,
  sink38,
  sink39,
  sink40,
  sink41,
  sink42,
  sink43,
  sink44,
  sink45,
  sink46,
  sink47,
  sink48,
  sink49,
  sink50,
  sink51,
  sink52,
  sink53,
  sink54,
  sink55,
  sink56,
  sink57,
  sink58,
  sink59,
  sink60,
  sink61,
  sink62,
  sink63,
  sink64,
  sink65,
  sink66,
  sink67,
  sink68,
  sink69,
  sink70,
  sink71,
  sink72,
  sink73,
  sink74,
  sink75,
  sink76,
  sink77,
  sink78,
  sink79,
  sink80,
  sink81,
  sink82,
  sink83,
  sink84,
  sink85,
  sink86,
  sink87,
  sink88,
  sink89,
  sink90,
  sink91,
  sink92,
  sink93,
  sink94,
  sink95,
  sink96,
  sink97,
  sink98,
  sink99,
  sink100,
  sink101,
  sink102,
  sink103,
  sink104,
  sink105,
  sink106,
  sink107,
  sink108,
  sink109,
  sink110,
  sink111,
  sink112,
  sink113,
  sink114,
  sink115,
  sink116,
  sink117,
  sink118,
  sink119,
  sink120,
  sink121,
  sink122,
  sink123,
  sink124,
  sink125,
  sink126,
  sink127,
  sink128,
  sink129,
  sink130,
  sink131,
  sink132,
  sink133,
  sink134,
  sink135,
  sink136,
  sink137,
  sink138,
  sink139,
  sink140,
  sink141,
  sink142,
  sink143,
  sink144,
  sink145,
  sink146,
  sink147,
  sink148,
  sink149,
  sink150,
  sink151,
  sink152,
  sink153,
  sink154,
  sink155,
  sink156,
  sink157,
  sink158,
  sink159,
  sink160,
  sink161,
  sink162,
  sink163,
  sink164,
  sink165,
  sink166,
  sink167,
  sink168,
  sink169,
  sink170,
  sink171,
  sink172,
  sink173,
  sink174,
  sink175,
  sink176,
  sink177,
  sink178,
  sink179,
  sink180,
  sink181,
  sink182,
  sink183,
  sink184,
  sink185,
  sink186,
  sink187,
  sink188,
  sink189,
  sink190,
  sink191,
  sink192,
  sink193,
  sink194,
  sink195,
  sink196,
  sink197,
  sink198,
  sink199,
  sink200,
  sink201,
  sink202,
  sink203,
  sink204,
  sink205,
  sink206,
  sink207,
  sink208,
  sink209,
  sink210,
  sink211,
  sink212,
  sink213,
  sink214,
  sink215,
  sink216,
  sink217,
  sink218,
  sink219,
  sink220,
  sink221,
  sink222,
  sink223,
  sink224,
  sink225,
  sink226,
  sink227,
  sink228,
  sink229,
  sink230,
  sink231,
  sink232,
  sink233,
  sink234,
  sink235,
  sink236,
  sink237,
  sink238,
  sink239,
  sink240,
  sink241,
  sink242,
  sink243,
  sink244,
  sink245,
  sink246,
  sink247,
  sink248,
  sink249,
  sink250,
  sink251,
  sink252,
  sink253,
  sink254,
  sink255,
  sink256,
  sink257,
  sink258,
  sink259,
  sink260,
  sink261,
  sink262,
  sink263,
  sink264,
  sink265,
  sink266
);
input clk;
output sink0;
output sink1;
output sink2;
output sink3;
output sink4;
output sink5;
output sink6;
output sink7;
output sink8;
output sink9;
output sink10;
output sink11;
output sink12;
output sink13;
output sink14;
output sink15;
output sink16;
output sink17;
output sink18;
output sink19;
output sink20;
output sink21;
output sink22;
output sink23;
output sink24;
output sink25;
output sink26;
output sink27;
output sink28;
output sink29;
output sink30;
output sink31;
output sink32;
output sink33;
output sink34;
output sink35;
output sink36;
output sink37;
output sink38;
output sink39;
output sink40;
output sink41;
output sink42;
output sink43;
output sink44;
output sink45;
output sink46;
output sink47;
output sink48;
output sink49;
output sink50;
output sink51;
output sink52;
output sink53;
output sink54;
output sink55;
output sink56;
output sink57;
output sink58;
output sink59;
output sink60;
output sink61;
output sink62;
output sink63;
output sink64;
output sink65;
output sink66;
output sink67;
output sink68;
output sink69;
output sink70;
output sink71;
output sink72;
output sink73;
output sink74;
output sink75;
output sink76;
output sink77;
output sink78;
output sink79;
output sink80;
output sink81;
output sink82;
output sink83;
output sink84;
output sink85;
output sink86;
output sink87;
output sink88;
output sink89;
output sink90;
output sink91;
output sink92;
output sink93;
output sink94;
output sink95;
output sink96;
output sink97;
output sink98;
output sink99;
output sink100;
output sink101;
output sink102;
output sink103;
output sink104;
output sink105;
output sink106;
output sink107;
output sink108;
output sink109;
output sink110;
output sink111;
output sink112;
output sink113;
output sink114;
output sink115;
output sink116;
output sink117;
output sink118;
output sink119;
output sink120;
output sink121;
output sink122;
output sink123;
output sink124;
output sink125;
output sink126;
output sink127;
output sink128;
output sink129;
output sink130;
output sink131;
output sink132;
output sink133;
output sink134;
output sink135;
output sink136;
output sink137;
output sink138;
output sink139;
output sink140;
output sink141;
output sink142;
output sink143;
output sink144;
output sink145;
output sink146;
output sink147;
output sink148;
output sink149;
output sink150;
output sink151;
output sink152;
output sink153;
output sink154;
output sink155;
output sink156;
output sink157;
output sink158;
output sink159;
output sink160;
output sink161;
output sink162;
output sink163;
output sink164;
output sink165;
output sink166;
output sink167;
output sink168;
output sink169;
output sink170;
output sink171;
output sink172;
output sink173;
output sink174;
output sink175;
output sink176;
output sink177;
output sink178;
output sink179;
output sink180;
output sink181;
output sink182;
output sink183;
output sink184;
output sink185;
output sink186;
output sink187;
output sink188;
output sink189;
output sink190;
output sink191;
output sink192;
output sink193;
output sink194;
output sink195;
output sink196;
output sink197;
output sink198;
output sink199;
output sink200;
output sink201;
output sink202;
output sink203;
output sink204;
output sink205;
output sink206;
output sink207;
output sink208;
output sink209;
output sink210;
output sink211;
output sink212;
output sink213;
output sink214;
output sink215;
output sink216;
output sink217;
output sink218;
output sink219;
output sink220;
output sink221;
output sink222;
output sink223;
output sink224;
output sink225;
output sink226;
output sink227;
output sink228;
output sink229;
output sink230;
output sink231;
output sink232;
output sink233;
output sink234;
output sink235;
output sink236;
output sink237;
output sink238;
output sink239;
output sink240;
output sink241;
output sink242;
output sink243;
output sink244;
output sink245;
output sink246;
output sink247;
output sink248;
output sink249;
output sink250;
output sink251;
output sink252;
output sink253;
output sink254;
output sink255;
output sink256;
output sink257;
output sink258;
output sink259;
output sink260;
output sink261;
output sink262;
output sink263;
output sink264;
output sink265;
output sink266;
  dff dff0 ( .clk(clk), .d(1'b0), .q(sink0));
  dff dff1 ( .clk(clk), .d(1'b0), .q(sink1));
  dff dff2 ( .clk(clk), .d(1'b0), .q(sink2));
  dff dff3 ( .clk(clk), .d(1'b0), .q(sink3));
  dff dff4 ( .clk(clk), .d(1'b0), .q(sink4));
  dff dff5 ( .clk(clk), .d(1'b0), .q(sink5));
  dff dff6 ( .clk(clk), .d(1'b0), .q(sink6));
  dff dff7 ( .clk(clk), .d(1'b0), .q(sink7));
  dff dff8 ( .clk(clk), .d(1'b0), .q(sink8));
  dff dff9 ( .clk(clk), .d(1'b0), .q(sink9));
  dff dff10 ( .clk(clk), .d(1'b0), .q(sink10));
  dff dff11 ( .clk(clk), .d(1'b0), .q(sink11));
  dff dff12 ( .clk(clk), .d(1'b0), .q(sink12));
  dff dff13 ( .clk(clk), .d(1'b0), .q(sink13));
  dff dff14 ( .clk(clk), .d(1'b0), .q(sink14));
  dff dff15 ( .clk(clk), .d(1'b0), .q(sink15));
  dff dff16 ( .clk(clk), .d(1'b0), .q(sink16));
  dff dff17 ( .clk(clk), .d(1'b0), .q(sink17));
  dff dff18 ( .clk(clk), .d(1'b0), .q(sink18));
  dff dff19 ( .clk(clk), .d(1'b0), .q(sink19));
  dff dff20 ( .clk(clk), .d(1'b0), .q(sink20));
  dff dff21 ( .clk(clk), .d(1'b0), .q(sink21));
  dff dff22 ( .clk(clk), .d(1'b0), .q(sink22));
  dff dff23 ( .clk(clk), .d(1'b0), .q(sink23));
  dff dff24 ( .clk(clk), .d(1'b0), .q(sink24));
  dff dff25 ( .clk(clk), .d(1'b0), .q(sink25));
  dff dff26 ( .clk(clk), .d(1'b0), .q(sink26));
  dff dff27 ( .clk(clk), .d(1'b0), .q(sink27));
  dff dff28 ( .clk(clk), .d(1'b0), .q(sink28));
  dff dff29 ( .clk(clk), .d(1'b0), .q(sink29));
  dff dff30 ( .clk(clk), .d(1'b0), .q(sink30));
  dff dff31 ( .clk(clk), .d(1'b0), .q(sink31));
  dff dff32 ( .clk(clk), .d(1'b0), .q(sink32));
  dff dff33 ( .clk(clk), .d(1'b0), .q(sink33));
  dff dff34 ( .clk(clk), .d(1'b0), .q(sink34));
  dff dff35 ( .clk(clk), .d(1'b0), .q(sink35));
  dff dff36 ( .clk(clk), .d(1'b0), .q(sink36));
  dff dff37 ( .clk(clk), .d(1'b0), .q(sink37));
  dff dff38 ( .clk(clk), .d(1'b0), .q(sink38));
  dff dff39 ( .clk(clk), .d(1'b0), .q(sink39));
  dff dff40 ( .clk(clk), .d(1'b0), .q(sink40));
  dff dff41 ( .clk(clk), .d(1'b0), .q(sink41));
  dff dff42 ( .clk(clk), .d(1'b0), .q(sink42));
  dff dff43 ( .clk(clk), .d(1'b0), .q(sink43));
  dff dff44 ( .clk(clk), .d(1'b0), .q(sink44));
  dff dff45 ( .clk(clk), .d(1'b0), .q(sink45));
  dff dff46 ( .clk(clk), .d(1'b0), .q(sink46));
  dff dff47 ( .clk(clk), .d(1'b0), .q(sink47));
  dff dff48 ( .clk(clk), .d(1'b0), .q(sink48));
  dff dff49 ( .clk(clk), .d(1'b0), .q(sink49));
  dff dff50 ( .clk(clk), .d(1'b0), .q(sink50));
  dff dff51 ( .clk(clk), .d(1'b0), .q(sink51));
  dff dff52 ( .clk(clk), .d(1'b0), .q(sink52));
  dff dff53 ( .clk(clk), .d(1'b0), .q(sink53));
  dff dff54 ( .clk(clk), .d(1'b0), .q(sink54));
  dff dff55 ( .clk(clk), .d(1'b0), .q(sink55));
  dff dff56 ( .clk(clk), .d(1'b0), .q(sink56));
  dff dff57 ( .clk(clk), .d(1'b0), .q(sink57));
  dff dff58 ( .clk(clk), .d(1'b0), .q(sink58));
  dff dff59 ( .clk(clk), .d(1'b0), .q(sink59));
  dff dff60 ( .clk(clk), .d(1'b0), .q(sink60));
  dff dff61 ( .clk(clk), .d(1'b0), .q(sink61));
  dff dff62 ( .clk(clk), .d(1'b0), .q(sink62));
  dff dff63 ( .clk(clk), .d(1'b0), .q(sink63));
  dff dff64 ( .clk(clk), .d(1'b0), .q(sink64));
  dff dff65 ( .clk(clk), .d(1'b0), .q(sink65));
  dff dff66 ( .clk(clk), .d(1'b0), .q(sink66));
  dff dff67 ( .clk(clk), .d(1'b0), .q(sink67));
  dff dff68 ( .clk(clk), .d(1'b0), .q(sink68));
  dff dff69 ( .clk(clk), .d(1'b0), .q(sink69));
  dff dff70 ( .clk(clk), .d(1'b0), .q(sink70));
  dff dff71 ( .clk(clk), .d(1'b0), .q(sink71));
  dff dff72 ( .clk(clk), .d(1'b0), .q(sink72));
  dff dff73 ( .clk(clk), .d(1'b0), .q(sink73));
  dff dff74 ( .clk(clk), .d(1'b0), .q(sink74));
  dff dff75 ( .clk(clk), .d(1'b0), .q(sink75));
  dff dff76 ( .clk(clk), .d(1'b0), .q(sink76));
  dff dff77 ( .clk(clk), .d(1'b0), .q(sink77));
  dff dff78 ( .clk(clk), .d(1'b0), .q(sink78));
  dff dff79 ( .clk(clk), .d(1'b0), .q(sink79));
  dff dff80 ( .clk(clk), .d(1'b0), .q(sink80));
  dff dff81 ( .clk(clk), .d(1'b0), .q(sink81));
  dff dff82 ( .clk(clk), .d(1'b0), .q(sink82));
  dff dff83 ( .clk(clk), .d(1'b0), .q(sink83));
  dff dff84 ( .clk(clk), .d(1'b0), .q(sink84));
  dff dff85 ( .clk(clk), .d(1'b0), .q(sink85));
  dff dff86 ( .clk(clk), .d(1'b0), .q(sink86));
  dff dff87 ( .clk(clk), .d(1'b0), .q(sink87));
  dff dff88 ( .clk(clk), .d(1'b0), .q(sink88));
  dff dff89 ( .clk(clk), .d(1'b0), .q(sink89));
  dff dff90 ( .clk(clk), .d(1'b0), .q(sink90));
  dff dff91 ( .clk(clk), .d(1'b0), .q(sink91));
  dff dff92 ( .clk(clk), .d(1'b0), .q(sink92));
  dff dff93 ( .clk(clk), .d(1'b0), .q(sink93));
  dff dff94 ( .clk(clk), .d(1'b0), .q(sink94));
  dff dff95 ( .clk(clk), .d(1'b0), .q(sink95));
  dff dff96 ( .clk(clk), .d(1'b0), .q(sink96));
  dff dff97 ( .clk(clk), .d(1'b0), .q(sink97));
  dff dff98 ( .clk(clk), .d(1'b0), .q(sink98));
  dff dff99 ( .clk(clk), .d(1'b0), .q(sink99));
  dff dff100 ( .clk(clk), .d(1'b0), .q(sink100));
  dff dff101 ( .clk(clk), .d(1'b0), .q(sink101));
  dff dff102 ( .clk(clk), .d(1'b0), .q(sink102));
  dff dff103 ( .clk(clk), .d(1'b0), .q(sink103));
  dff dff104 ( .clk(clk), .d(1'b0), .q(sink104));
  dff dff105 ( .clk(clk), .d(1'b0), .q(sink105));
  dff dff106 ( .clk(clk), .d(1'b0), .q(sink106));
  dff dff107 ( .clk(clk), .d(1'b0), .q(sink107));
  dff dff108 ( .clk(clk), .d(1'b0), .q(sink108));
  dff dff109 ( .clk(clk), .d(1'b0), .q(sink109));
  dff dff110 ( .clk(clk), .d(1'b0), .q(sink110));
  dff dff111 ( .clk(clk), .d(1'b0), .q(sink111));
  dff dff112 ( .clk(clk), .d(1'b0), .q(sink112));
  dff dff113 ( .clk(clk), .d(1'b0), .q(sink113));
  dff dff114 ( .clk(clk), .d(1'b0), .q(sink114));
  dff dff115 ( .clk(clk), .d(1'b0), .q(sink115));
  dff dff116 ( .clk(clk), .d(1'b0), .q(sink116));
  dff dff117 ( .clk(clk), .d(1'b0), .q(sink117));
  dff dff118 ( .clk(clk), .d(1'b0), .q(sink118));
  dff dff119 ( .clk(clk), .d(1'b0), .q(sink119));
  dff dff120 ( .clk(clk), .d(1'b0), .q(sink120));
  dff dff121 ( .clk(clk), .d(1'b0), .q(sink121));
  dff dff122 ( .clk(clk), .d(1'b0), .q(sink122));
  dff dff123 ( .clk(clk), .d(1'b0), .q(sink123));
  dff dff124 ( .clk(clk), .d(1'b0), .q(sink124));
  dff dff125 ( .clk(clk), .d(1'b0), .q(sink125));
  dff dff126 ( .clk(clk), .d(1'b0), .q(sink126));
  dff dff127 ( .clk(clk), .d(1'b0), .q(sink127));
  dff dff128 ( .clk(clk), .d(1'b0), .q(sink128));
  dff dff129 ( .clk(clk), .d(1'b0), .q(sink129));
  dff dff130 ( .clk(clk), .d(1'b0), .q(sink130));
  dff dff131 ( .clk(clk), .d(1'b0), .q(sink131));
  dff dff132 ( .clk(clk), .d(1'b0), .q(sink132));
  dff dff133 ( .clk(clk), .d(1'b0), .q(sink133));
  dff dff134 ( .clk(clk), .d(1'b0), .q(sink134));
  dff dff135 ( .clk(clk), .d(1'b0), .q(sink135));
  dff dff136 ( .clk(clk), .d(1'b0), .q(sink136));
  dff dff137 ( .clk(clk), .d(1'b0), .q(sink137));
  dff dff138 ( .clk(clk), .d(1'b0), .q(sink138));
  dff dff139 ( .clk(clk), .d(1'b0), .q(sink139));
  dff dff140 ( .clk(clk), .d(1'b0), .q(sink140));
  dff dff141 ( .clk(clk), .d(1'b0), .q(sink141));
  dff dff142 ( .clk(clk), .d(1'b0), .q(sink142));
  dff dff143 ( .clk(clk), .d(1'b0), .q(sink143));
  dff dff144 ( .clk(clk), .d(1'b0), .q(sink144));
  dff dff145 ( .clk(clk), .d(1'b0), .q(sink145));
  dff dff146 ( .clk(clk), .d(1'b0), .q(sink146));
  dff dff147 ( .clk(clk), .d(1'b0), .q(sink147));
  dff dff148 ( .clk(clk), .d(1'b0), .q(sink148));
  dff dff149 ( .clk(clk), .d(1'b0), .q(sink149));
  dff dff150 ( .clk(clk), .d(1'b0), .q(sink150));
  dff dff151 ( .clk(clk), .d(1'b0), .q(sink151));
  dff dff152 ( .clk(clk), .d(1'b0), .q(sink152));
  dff dff153 ( .clk(clk), .d(1'b0), .q(sink153));
  dff dff154 ( .clk(clk), .d(1'b0), .q(sink154));
  dff dff155 ( .clk(clk), .d(1'b0), .q(sink155));
  dff dff156 ( .clk(clk), .d(1'b0), .q(sink156));
  dff dff157 ( .clk(clk), .d(1'b0), .q(sink157));
  dff dff158 ( .clk(clk), .d(1'b0), .q(sink158));
  dff dff159 ( .clk(clk), .d(1'b0), .q(sink159));
  dff dff160 ( .clk(clk), .d(1'b0), .q(sink160));
  dff dff161 ( .clk(clk), .d(1'b0), .q(sink161));
  dff dff162 ( .clk(clk), .d(1'b0), .q(sink162));
  dff dff163 ( .clk(clk), .d(1'b0), .q(sink163));
  dff dff164 ( .clk(clk), .d(1'b0), .q(sink164));
  dff dff165 ( .clk(clk), .d(1'b0), .q(sink165));
  dff dff166 ( .clk(clk), .d(1'b0), .q(sink166));
  dff dff167 ( .clk(clk), .d(1'b0), .q(sink167));
  dff dff168 ( .clk(clk), .d(1'b0), .q(sink168));
  dff dff169 ( .clk(clk), .d(1'b0), .q(sink169));
  dff dff170 ( .clk(clk), .d(1'b0), .q(sink170));
  dff dff171 ( .clk(clk), .d(1'b0), .q(sink171));
  dff dff172 ( .clk(clk), .d(1'b0), .q(sink172));
  dff dff173 ( .clk(clk), .d(1'b0), .q(sink173));
  dff dff174 ( .clk(clk), .d(1'b0), .q(sink174));
  dff dff175 ( .clk(clk), .d(1'b0), .q(sink175));
  dff dff176 ( .clk(clk), .d(1'b0), .q(sink176));
  dff dff177 ( .clk(clk), .d(1'b0), .q(sink177));
  dff dff178 ( .clk(clk), .d(1'b0), .q(sink178));
  dff dff179 ( .clk(clk), .d(1'b0), .q(sink179));
  dff dff180 ( .clk(clk), .d(1'b0), .q(sink180));
  dff dff181 ( .clk(clk), .d(1'b0), .q(sink181));
  dff dff182 ( .clk(clk), .d(1'b0), .q(sink182));
  dff dff183 ( .clk(clk), .d(1'b0), .q(sink183));
  dff dff184 ( .clk(clk), .d(1'b0), .q(sink184));
  dff dff185 ( .clk(clk), .d(1'b0), .q(sink185));
  dff dff186 ( .clk(clk), .d(1'b0), .q(sink186));
  dff dff187 ( .clk(clk), .d(1'b0), .q(sink187));
  dff dff188 ( .clk(clk), .d(1'b0), .q(sink188));
  dff dff189 ( .clk(clk), .d(1'b0), .q(sink189));
  dff dff190 ( .clk(clk), .d(1'b0), .q(sink190));
  dff dff191 ( .clk(clk), .d(1'b0), .q(sink191));
  dff dff192 ( .clk(clk), .d(1'b0), .q(sink192));
  dff dff193 ( .clk(clk), .d(1'b0), .q(sink193));
  dff dff194 ( .clk(clk), .d(1'b0), .q(sink194));
  dff dff195 ( .clk(clk), .d(1'b0), .q(sink195));
  dff dff196 ( .clk(clk), .d(1'b0), .q(sink196));
  dff dff197 ( .clk(clk), .d(1'b0), .q(sink197));
  dff dff198 ( .clk(clk), .d(1'b0), .q(sink198));
  dff dff199 ( .clk(clk), .d(1'b0), .q(sink199));
  dff dff200 ( .clk(clk), .d(1'b0), .q(sink200));
  dff dff201 ( .clk(clk), .d(1'b0), .q(sink201));
  dff dff202 ( .clk(clk), .d(1'b0), .q(sink202));
  dff dff203 ( .clk(clk), .d(1'b0), .q(sink203));
  dff dff204 ( .clk(clk), .d(1'b0), .q(sink204));
  dff dff205 ( .clk(clk), .d(1'b0), .q(sink205));
  dff dff206 ( .clk(clk), .d(1'b0), .q(sink206));
  dff dff207 ( .clk(clk), .d(1'b0), .q(sink207));
  dff dff208 ( .clk(clk), .d(1'b0), .q(sink208));
  dff dff209 ( .clk(clk), .d(1'b0), .q(sink209));
  dff dff210 ( .clk(clk), .d(1'b0), .q(sink210));
  dff dff211 ( .clk(clk), .d(1'b0), .q(sink211));
  dff dff212 ( .clk(clk), .d(1'b0), .q(sink212));
  dff dff213 ( .clk(clk), .d(1'b0), .q(sink213));
  dff dff214 ( .clk(clk), .d(1'b0), .q(sink214));
  dff dff215 ( .clk(clk), .d(1'b0), .q(sink215));
  dff dff216 ( .clk(clk), .d(1'b0), .q(sink216));
  dff dff217 ( .clk(clk), .d(1'b0), .q(sink217));
  dff dff218 ( .clk(clk), .d(1'b0), .q(sink218));
  dff dff219 ( .clk(clk), .d(1'b0), .q(sink219));
  dff dff220 ( .clk(clk), .d(1'b0), .q(sink220));
  dff dff221 ( .clk(clk), .d(1'b0), .q(sink221));
  dff dff222 ( .clk(clk), .d(1'b0), .q(sink222));
  dff dff223 ( .clk(clk), .d(1'b0), .q(sink223));
  dff dff224 ( .clk(clk), .d(1'b0), .q(sink224));
  dff dff225 ( .clk(clk), .d(1'b0), .q(sink225));
  dff dff226 ( .clk(clk), .d(1'b0), .q(sink226));
  dff dff227 ( .clk(clk), .d(1'b0), .q(sink227));
  dff dff228 ( .clk(clk), .d(1'b0), .q(sink228));
  dff dff229 ( .clk(clk), .d(1'b0), .q(sink229));
  dff dff230 ( .clk(clk), .d(1'b0), .q(sink230));
  dff dff231 ( .clk(clk), .d(1'b0), .q(sink231));
  dff dff232 ( .clk(clk), .d(1'b0), .q(sink232));
  dff dff233 ( .clk(clk), .d(1'b0), .q(sink233));
  dff dff234 ( .clk(clk), .d(1'b0), .q(sink234));
  dff dff235 ( .clk(clk), .d(1'b0), .q(sink235));
  dff dff236 ( .clk(clk), .d(1'b0), .q(sink236));
  dff dff237 ( .clk(clk), .d(1'b0), .q(sink237));
  dff dff238 ( .clk(clk), .d(1'b0), .q(sink238));
  dff dff239 ( .clk(clk), .d(1'b0), .q(sink239));
  dff dff240 ( .clk(clk), .d(1'b0), .q(sink240));
  dff dff241 ( .clk(clk), .d(1'b0), .q(sink241));
  dff dff242 ( .clk(clk), .d(1'b0), .q(sink242));
  dff dff243 ( .clk(clk), .d(1'b0), .q(sink243));
  dff dff244 ( .clk(clk), .d(1'b0), .q(sink244));
  dff dff245 ( .clk(clk), .d(1'b0), .q(sink245));
  dff dff246 ( .clk(clk), .d(1'b0), .q(sink246));
  dff dff247 ( .clk(clk), .d(1'b0), .q(sink247));
  dff dff248 ( .clk(clk), .d(1'b0), .q(sink248));
  dff dff249 ( .clk(clk), .d(1'b0), .q(sink249));
  dff dff250 ( .clk(clk), .d(1'b0), .q(sink250));
  dff dff251 ( .clk(clk), .d(1'b0), .q(sink251));
  dff dff252 ( .clk(clk), .d(1'b0), .q(sink252));
  dff dff253 ( .clk(clk), .d(1'b0), .q(sink253));
  dff dff254 ( .clk(clk), .d(1'b0), .q(sink254));
  dff dff255 ( .clk(clk), .d(1'b0), .q(sink255));
  dff dff256 ( .clk(clk), .d(1'b0), .q(sink256));
  dff dff257 ( .clk(clk), .d(1'b0), .q(sink257));
  dff dff258 ( .clk(clk), .d(1'b0), .q(sink258));
  dff dff259 ( .clk(clk), .d(1'b0), .q(sink259));
  dff dff260 ( .clk(clk), .d(1'b0), .q(sink260));
  dff dff261 ( .clk(clk), .d(1'b0), .q(sink261));
  dff dff262 ( .clk(clk), .d(1'b0), .q(sink262));
  dff dff263 ( .clk(clk), .d(1'b0), .q(sink263));
  dff dff264 ( .clk(clk), .d(1'b0), .q(sink264));
  dff dff265 ( .clk(clk), .d(1'b0), .q(sink265));
  dff dff266 ( .clk(clk), .d(1'b0), .q(sink266));
endmodule