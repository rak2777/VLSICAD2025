module top (input clk);
  DFF u_ff_0.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_1.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_2.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_3.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_4.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_5.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_6.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_7.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_8.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_9.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_10.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_11.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_12.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_13.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_14.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_15.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_16.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_17.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_18.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_19.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_20.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_21.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_22.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_23.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_24.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_25.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_26.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_27.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_28.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_29.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_30.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_31.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_32.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_33.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_34.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_35.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_36.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_37.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_38.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_39.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_40.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_41.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_42.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_43.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_44.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_45.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_46.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_47.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_48.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_49.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_50.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_51.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_52.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_53.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_54.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_55.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_56.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_57.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_58.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_59.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_60.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_61.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_62.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_63.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_64.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_65.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_66.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_67.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_68.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_69.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_70.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_71.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_72.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_73.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_74.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_75.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_76.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_77.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_78.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_79.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_80.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_81.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_82.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_83.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_84.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_85.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_86.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_87.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_88.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_89.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_90.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_91.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_92.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_93.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_94.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_95.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_96.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_97.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_98.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_99.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_100.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_101.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_102.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_103.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_104.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_105.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_106.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_107.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_108.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_109.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_110.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_111.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_112.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_113.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_114.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_115.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_116.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_117.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_118.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_119.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_120.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_121.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_122.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_123.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_124.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_125.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_126.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_127.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_128.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_129.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_130.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_131.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_132.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_133.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_134.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_135.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_136.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_137.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_138.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_139.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_140.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_141.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_142.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_143.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_144.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_145.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_146.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_147.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_148.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_149.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_150.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_151.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_152.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_153.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_154.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_155.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_156.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_157.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_158.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_159.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_160.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_161.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_162.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_163.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_164.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_165.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_166.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_167.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_168.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_169.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_170.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_171.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_172.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_173.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_174.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_175.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_176.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_177.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_178.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_179.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_180.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_181.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_182.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_183.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_184.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_185.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_186.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_187.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_188.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_189.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_190.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_191.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_192.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_193.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_194.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_195.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_196.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_197.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_198.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_199.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_200.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_201.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_202.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_203.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_204.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_205.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_206.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_207.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_208.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_209.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_210.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_211.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_212.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_213.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_214.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_215.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_216.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_217.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_218.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_219.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_220.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_221.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_222.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_223.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_224.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_225.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_226.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_227.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_228.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_229.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_230.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_231.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_232.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_233.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_234.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_235.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_236.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_237.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_238.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_239.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_240.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_241.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_242.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_243.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_244.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_245.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_246.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_247.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_248.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_249.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_250.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_251.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_252.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_253.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_254.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_255.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_256.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_257.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_258.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_259.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_260.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_261.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_262.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_263.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_264.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_265.0 (.clk(clk), .d(1'b0), .q());
  DFF u_ff_266.0 (.clk(clk), .d(1'b0), .q());
endmodule