module clock_tree (
    clk,
    out_0, 
    out_1, 
    out_2, 
    out_3, 
    out_4, 
    out_5, 
    out_6, 
    out_7, 
    out_8, 
    out_9, 
    out_10, 
    out_11, 
    out_12, 
    out_13, 
    out_14, 
    out_15, 
    out_16, 
    out_17, 
    out_18, 
    out_19, 
    out_20, 
    out_21, 
    out_22, 
    out_23, 
    out_24, 
    out_25, 
    out_26, 
    out_27, 
    out_28, 
    out_29, 
    out_30, 
    out_31, 
    out_32, 
    out_33, 
    out_34, 
    out_35, 
    out_36, 
    out_37, 
    out_38, 
    out_39, 
    out_40, 
    out_41, 
    out_42, 
    out_43, 
    out_44, 
    out_45, 
    out_46, 
    out_47, 
    out_48, 
    out_49, 
    out_50, 
    out_51, 
    out_52, 
    out_53, 
    out_54, 
    out_55, 
    out_56, 
    out_57, 
    out_58, 
    out_59, 
    out_60, 
    out_61, 
    out_62, 
    out_63, 
    out_64, 
    out_65, 
    out_66, 
    out_67, 
    out_68, 
    out_69, 
    out_70, 
    out_71, 
    out_72, 
    out_73, 
    out_74, 
    out_75, 
    out_76, 
    out_77, 
    out_78, 
    out_79, 
    out_80, 
    out_81, 
    out_82, 
    out_83, 
    out_84, 
    out_85, 
    out_86, 
    out_87, 
    out_88, 
    out_89, 
    out_90, 
    out_91, 
    out_92, 
    out_93, 
    out_94, 
    out_95, 
    out_96, 
    out_97, 
    out_98, 
    out_99, 
    out_100, 
    out_101, 
    out_102, 
    out_103, 
    out_104, 
    out_105, 
    out_106, 
    out_107, 
    out_108, 
    out_109, 
    out_110, 
    out_111, 
    out_112, 
    out_113, 
    out_114, 
    out_115, 
    out_116, 
    out_117, 
    out_118, 
    out_119, 
    out_120, 
    out_121, 
    out_122, 
    out_123, 
    out_124, 
    out_125, 
    out_126, 
    out_127, 
    out_128, 
    out_129, 
    out_130, 
    out_131, 
    out_132, 
    out_133, 
    out_134, 
    out_135, 
    out_136, 
    out_137, 
    out_138, 
    out_139, 
    out_140, 
    out_141, 
    out_142, 
    out_143, 
    out_144, 
    out_145, 
    out_146, 
    out_147, 
    out_148, 
    out_149, 
    out_150, 
    out_151, 
    out_152, 
    out_153, 
    out_154, 
    out_155, 
    out_156, 
    out_157, 
    out_158, 
    out_159, 
    out_160, 
    out_161, 
    out_162, 
    out_163, 
    out_164, 
    out_165, 
    out_166, 
    out_167, 
    out_168, 
    out_169, 
    out_170, 
    out_171, 
    out_172, 
    out_173, 
    out_174, 
    out_175, 
    out_176, 
    out_177, 
    out_178, 
    out_179, 
    out_180, 
    out_181, 
    out_182, 
    out_183, 
    out_184, 
    out_185, 
    out_186, 
    out_187, 
    out_188, 
    out_189, 
    out_190, 
    out_191, 
    out_192, 
    out_193, 
    out_194, 
    out_195, 
    out_196, 
    out_197, 
    out_198, 
    out_199, 
    out_200, 
    out_201, 
    out_202, 
    out_203, 
    out_204, 
    out_205, 
    out_206, 
    out_207, 
    out_208, 
    out_209, 
    out_210, 
    out_211, 
    out_212, 
    out_213, 
    out_214, 
    out_215, 
    out_216, 
    out_217, 
    out_218, 
    out_219, 
    out_220, 
    out_221, 
    out_222, 
    out_223, 
    out_224, 
    out_225, 
    out_226, 
    out_227, 
    out_228, 
    out_229, 
    out_230, 
    out_231, 
    out_232, 
    out_233, 
    out_234, 
    out_235, 
    out_236, 
    out_237, 
    out_238, 
    out_239, 
    out_240, 
    out_241, 
    out_242, 
    out_243, 
    out_244, 
    out_245, 
    out_246, 
    out_247, 
    out_248, 
    out_249, 
    out_250, 
    out_251, 
    out_252, 
    out_253, 
    out_254, 
    out_255, 
    out_256, 
    out_257, 
    out_258, 
    out_259, 
    out_260, 
    out_261, 
    out_262, 
    out_263, 
    out_264, 
    out_265, 
    out_266, 
);

input clk;
output out_0;
output out_1;
output out_2;
output out_3;
output out_4;
output out_5;
output out_6;
output out_7;
output out_8;
output out_9;
output out_10;
output out_11;
output out_12;
output out_13;
output out_14;
output out_15;
output out_16;
output out_17;
output out_18;
output out_19;
output out_20;
output out_21;
output out_22;
output out_23;
output out_24;
output out_25;
output out_26;
output out_27;
output out_28;
output out_29;
output out_30;
output out_31;
output out_32;
output out_33;
output out_34;
output out_35;
output out_36;
output out_37;
output out_38;
output out_39;
output out_40;
output out_41;
output out_42;
output out_43;
output out_44;
output out_45;
output out_46;
output out_47;
output out_48;
output out_49;
output out_50;
output out_51;
output out_52;
output out_53;
output out_54;
output out_55;
output out_56;
output out_57;
output out_58;
output out_59;
output out_60;
output out_61;
output out_62;
output out_63;
output out_64;
output out_65;
output out_66;
output out_67;
output out_68;
output out_69;
output out_70;
output out_71;
output out_72;
output out_73;
output out_74;
output out_75;
output out_76;
output out_77;
output out_78;
output out_79;
output out_80;
output out_81;
output out_82;
output out_83;
output out_84;
output out_85;
output out_86;
output out_87;
output out_88;
output out_89;
output out_90;
output out_91;
output out_92;
output out_93;
output out_94;
output out_95;
output out_96;
output out_97;
output out_98;
output out_99;
output out_100;
output out_101;
output out_102;
output out_103;
output out_104;
output out_105;
output out_106;
output out_107;
output out_108;
output out_109;
output out_110;
output out_111;
output out_112;
output out_113;
output out_114;
output out_115;
output out_116;
output out_117;
output out_118;
output out_119;
output out_120;
output out_121;
output out_122;
output out_123;
output out_124;
output out_125;
output out_126;
output out_127;
output out_128;
output out_129;
output out_130;
output out_131;
output out_132;
output out_133;
output out_134;
output out_135;
output out_136;
output out_137;
output out_138;
output out_139;
output out_140;
output out_141;
output out_142;
output out_143;
output out_144;
output out_145;
output out_146;
output out_147;
output out_148;
output out_149;
output out_150;
output out_151;
output out_152;
output out_153;
output out_154;
output out_155;
output out_156;
output out_157;
output out_158;
output out_159;
output out_160;
output out_161;
output out_162;
output out_163;
output out_164;
output out_165;
output out_166;
output out_167;
output out_168;
output out_169;
output out_170;
output out_171;
output out_172;
output out_173;
output out_174;
output out_175;
output out_176;
output out_177;
output out_178;
output out_179;
output out_180;
output out_181;
output out_182;
output out_183;
output out_184;
output out_185;
output out_186;
output out_187;
output out_188;
output out_189;
output out_190;
output out_191;
output out_192;
output out_193;
output out_194;
output out_195;
output out_196;
output out_197;
output out_198;
output out_199;
output out_200;
output out_201;
output out_202;
output out_203;
output out_204;
output out_205;
output out_206;
output out_207;
output out_208;
output out_209;
output out_210;
output out_211;
output out_212;
output out_213;
output out_214;
output out_215;
output out_216;
output out_217;
output out_218;
output out_219;
output out_220;
output out_221;
output out_222;
output out_223;
output out_224;
output out_225;
output out_226;
output out_227;
output out_228;
output out_229;
output out_230;
output out_231;
output out_232;
output out_233;
output out_234;
output out_235;
output out_236;
output out_237;
output out_238;
output out_239;
output out_240;
output out_241;
output out_242;
output out_243;
output out_244;
output out_245;
output out_246;
output out_247;
output out_248;
output out_249;
output out_250;
output out_251;
output out_252;
output out_253;
output out_254;
output out_255;
output out_256;
output out_257;
output out_258;
output out_259;
output out_260;
output out_261;
output out_262;
output out_263;
output out_264;
output out_265;
output out_266;

nand2x1 I1 ( .B(out_0), .A(out_1), .Z(net_1) );
nand2x1 I2 ( .B(out_0), .A(out_2), .Z(net_2) );
nand2x1 I3 ( .B(out_1), .A(out_3), .Z(net_3) );
nand2x1 I4 ( .B(out_1), .A(out_4), .Z(net_4) );
nand2x1 I5 ( .B(out_2), .A(out_5), .Z(net_5) );
nand2x1 I6 ( .B(out_2), .A(out_6), .Z(net_6) );
nand2x1 I7 ( .B(out_3), .A(out_7), .Z(net_7) );
nand2x1 I8 ( .B(out_3), .A(out_8), .Z(net_8) );
nand2x1 I9 ( .B(out_4), .A(out_9), .Z(net_9) );
nand2x1 I10 ( .B(out_4), .A(out_10), .Z(net_10) );
nand2x1 I11 ( .B(out_5), .A(out_11), .Z(net_11) );
nand2x1 I12 ( .B(out_5), .A(out_12), .Z(net_12) );
nand2x1 I13 ( .B(out_6), .A(out_13), .Z(net_13) );
nand2x1 I14 ( .B(out_6), .A(out_14), .Z(net_14) );
nand2x1 I15 ( .B(out_7), .A(out_15), .Z(net_15) );
nand2x1 I16 ( .B(out_7), .A(out_16), .Z(net_16) );
nand2x1 I17 ( .B(out_8), .A(out_17), .Z(net_17) );
nand2x1 I18 ( .B(out_8), .A(out_18), .Z(net_18) );
nand2x1 I19 ( .B(out_9), .A(out_19), .Z(net_19) );
nand2x1 I20 ( .B(out_9), .A(out_20), .Z(net_20) );
nand2x1 I21 ( .B(out_10), .A(out_21), .Z(net_21) );
nand2x1 I22 ( .B(out_10), .A(out_22), .Z(net_22) );
nand2x1 I23 ( .B(out_11), .A(out_23), .Z(net_23) );
nand2x1 I24 ( .B(out_11), .A(out_24), .Z(net_24) );
nand2x1 I25 ( .B(out_12), .A(out_25), .Z(net_25) );
nand2x1 I26 ( .B(out_12), .A(out_26), .Z(net_26) );
nand2x1 I27 ( .B(out_13), .A(out_27), .Z(net_27) );
nand2x1 I28 ( .B(out_13), .A(out_28), .Z(net_28) );
nand2x1 I29 ( .B(out_14), .A(out_29), .Z(net_29) );
nand2x1 I30 ( .B(out_14), .A(out_30), .Z(net_30) );
nand2x1 I31 ( .B(out_15), .A(out_31), .Z(net_31) );
nand2x1 I32 ( .B(out_15), .A(out_32), .Z(net_32) );
nand2x1 I33 ( .B(out_16), .A(out_33), .Z(net_33) );
nand2x1 I34 ( .B(out_16), .A(out_34), .Z(net_34) );
nand2x1 I35 ( .B(out_17), .A(out_35), .Z(net_35) );
nand2x1 I36 ( .B(out_17), .A(out_36), .Z(net_36) );
nand2x1 I37 ( .B(out_18), .A(out_37), .Z(net_37) );
nand2x1 I38 ( .B(out_18), .A(out_38), .Z(net_38) );
nand2x1 I39 ( .B(out_19), .A(out_39), .Z(net_39) );
nand2x1 I40 ( .B(out_19), .A(out_40), .Z(net_40) );
nand2x1 I41 ( .B(out_20), .A(out_41), .Z(net_41) );
nand2x1 I42 ( .B(out_20), .A(out_42), .Z(net_42) );
nand2x1 I43 ( .B(out_21), .A(out_43), .Z(net_43) );
nand2x1 I44 ( .B(out_21), .A(out_44), .Z(net_44) );
nand2x1 I45 ( .B(out_22), .A(out_45), .Z(net_45) );
nand2x1 I46 ( .B(out_22), .A(out_46), .Z(net_46) );
nand2x1 I47 ( .B(out_23), .A(out_47), .Z(net_47) );
nand2x1 I48 ( .B(out_23), .A(out_48), .Z(net_48) );
nand2x1 I49 ( .B(out_24), .A(out_49), .Z(net_49) );
nand2x1 I50 ( .B(out_24), .A(out_50), .Z(net_50) );
nand2x1 I51 ( .B(out_25), .A(out_51), .Z(net_51) );
nand2x1 I52 ( .B(out_25), .A(out_52), .Z(net_52) );
nand2x1 I53 ( .B(out_26), .A(out_53), .Z(net_53) );
nand2x1 I54 ( .B(out_26), .A(out_54), .Z(net_54) );
nand2x1 I55 ( .B(out_27), .A(out_55), .Z(net_55) );
nand2x1 I56 ( .B(out_27), .A(out_56), .Z(net_56) );
nand2x1 I57 ( .B(out_28), .A(out_57), .Z(net_57) );
nand2x1 I58 ( .B(out_28), .A(out_58), .Z(net_58) );
nand2x1 I59 ( .B(out_29), .A(out_59), .Z(net_59) );
nand2x1 I60 ( .B(out_29), .A(out_60), .Z(net_60) );
nand2x1 I61 ( .B(out_30), .A(out_61), .Z(net_61) );
nand2x1 I62 ( .B(out_30), .A(out_62), .Z(net_62) );
nand2x1 I63 ( .B(out_31), .A(out_63), .Z(net_63) );
nand2x1 I64 ( .B(out_31), .A(out_64), .Z(net_64) );
nand2x1 I65 ( .B(out_32), .A(out_65), .Z(net_65) );
nand2x1 I66 ( .B(out_32), .A(out_66), .Z(net_66) );
nand2x1 I67 ( .B(out_33), .A(out_67), .Z(net_67) );
nand2x1 I68 ( .B(out_33), .A(out_68), .Z(net_68) );
nand2x1 I69 ( .B(out_34), .A(out_69), .Z(net_69) );
nand2x1 I70 ( .B(out_34), .A(out_70), .Z(net_70) );
nand2x1 I71 ( .B(out_35), .A(out_71), .Z(net_71) );
nand2x1 I72 ( .B(out_35), .A(out_72), .Z(net_72) );
nand2x1 I73 ( .B(out_36), .A(out_73), .Z(net_73) );
nand2x1 I74 ( .B(out_36), .A(out_74), .Z(net_74) );
nand2x1 I75 ( .B(out_37), .A(out_75), .Z(net_75) );
nand2x1 I76 ( .B(out_37), .A(out_76), .Z(net_76) );
nand2x1 I77 ( .B(out_38), .A(out_77), .Z(net_77) );
nand2x1 I78 ( .B(out_38), .A(out_78), .Z(net_78) );
nand2x1 I79 ( .B(out_39), .A(out_79), .Z(net_79) );
nand2x1 I80 ( .B(out_39), .A(out_80), .Z(net_80) );
nand2x1 I81 ( .B(out_40), .A(out_81), .Z(net_81) );
nand2x1 I82 ( .B(out_40), .A(out_82), .Z(net_82) );
nand2x1 I83 ( .B(out_41), .A(out_83), .Z(net_83) );
nand2x1 I84 ( .B(out_41), .A(out_84), .Z(net_84) );
nand2x1 I85 ( .B(out_42), .A(out_85), .Z(net_85) );
nand2x1 I86 ( .B(out_42), .A(out_86), .Z(net_86) );
nand2x1 I87 ( .B(out_43), .A(out_87), .Z(net_87) );
nand2x1 I88 ( .B(out_43), .A(out_88), .Z(net_88) );
nand2x1 I89 ( .B(out_44), .A(out_89), .Z(net_89) );
nand2x1 I90 ( .B(out_44), .A(out_90), .Z(net_90) );
nand2x1 I91 ( .B(out_45), .A(out_91), .Z(net_91) );
nand2x1 I92 ( .B(out_45), .A(out_92), .Z(net_92) );
nand2x1 I93 ( .B(out_46), .A(out_93), .Z(net_93) );
nand2x1 I94 ( .B(out_46), .A(out_94), .Z(net_94) );
nand2x1 I95 ( .B(out_47), .A(out_95), .Z(net_95) );
nand2x1 I96 ( .B(out_47), .A(out_96), .Z(net_96) );
nand2x1 I97 ( .B(out_48), .A(out_97), .Z(net_97) );
nand2x1 I98 ( .B(out_48), .A(out_98), .Z(net_98) );
nand2x1 I99 ( .B(out_49), .A(out_99), .Z(net_99) );
nand2x1 I100 ( .B(out_49), .A(out_100), .Z(net_100) );
nand2x1 I101 ( .B(out_50), .A(out_101), .Z(net_101) );
nand2x1 I102 ( .B(out_50), .A(out_102), .Z(net_102) );
nand2x1 I103 ( .B(out_51), .A(out_103), .Z(net_103) );
nand2x1 I104 ( .B(out_51), .A(out_104), .Z(net_104) );
nand2x1 I105 ( .B(out_52), .A(out_105), .Z(net_105) );
nand2x1 I106 ( .B(out_52), .A(out_106), .Z(net_106) );
nand2x1 I107 ( .B(out_53), .A(out_107), .Z(net_107) );
nand2x1 I108 ( .B(out_53), .A(out_108), .Z(net_108) );
nand2x1 I109 ( .B(out_54), .A(out_109), .Z(net_109) );
nand2x1 I110 ( .B(out_54), .A(out_110), .Z(net_110) );
nand2x1 I111 ( .B(out_55), .A(out_111), .Z(net_111) );
nand2x1 I112 ( .B(out_55), .A(out_112), .Z(net_112) );
nand2x1 I113 ( .B(out_56), .A(out_113), .Z(net_113) );
nand2x1 I114 ( .B(out_56), .A(out_114), .Z(net_114) );
nand2x1 I115 ( .B(out_57), .A(out_115), .Z(net_115) );
nand2x1 I116 ( .B(out_57), .A(out_116), .Z(net_116) );
nand2x1 I117 ( .B(out_58), .A(out_117), .Z(net_117) );
nand2x1 I118 ( .B(out_58), .A(out_118), .Z(net_118) );
nand2x1 I119 ( .B(out_59), .A(out_119), .Z(net_119) );
nand2x1 I120 ( .B(out_59), .A(out_120), .Z(net_120) );
nand2x1 I121 ( .B(out_60), .A(out_121), .Z(net_121) );
nand2x1 I122 ( .B(out_60), .A(out_122), .Z(net_122) );
nand2x1 I123 ( .B(out_61), .A(out_123), .Z(net_123) );
nand2x1 I124 ( .B(out_61), .A(out_124), .Z(net_124) );
nand2x1 I125 ( .B(out_62), .A(out_125), .Z(net_125) );
nand2x1 I126 ( .B(out_62), .A(out_126), .Z(net_126) );
nand2x1 I127 ( .B(out_63), .A(out_127), .Z(net_127) );
nand2x1 I128 ( .B(out_63), .A(out_128), .Z(net_128) );
nand2x1 I129 ( .B(out_64), .A(out_129), .Z(net_129) );
nand2x1 I130 ( .B(out_64), .A(out_130), .Z(net_130) );
nand2x1 I131 ( .B(out_65), .A(out_131), .Z(net_131) );
nand2x1 I132 ( .B(out_65), .A(out_132), .Z(net_132) );
nand2x1 I133 ( .B(out_66), .A(out_133), .Z(net_133) );
nand2x1 I134 ( .B(out_66), .A(out_134), .Z(net_134) );
nand2x1 I135 ( .B(out_67), .A(out_135), .Z(net_135) );
nand2x1 I136 ( .B(out_67), .A(out_136), .Z(net_136) );
nand2x1 I137 ( .B(out_68), .A(out_137), .Z(net_137) );
nand2x1 I138 ( .B(out_68), .A(out_138), .Z(net_138) );
nand2x1 I139 ( .B(out_69), .A(out_139), .Z(net_139) );
nand2x1 I140 ( .B(out_69), .A(out_140), .Z(net_140) );
nand2x1 I141 ( .B(out_70), .A(out_141), .Z(net_141) );
nand2x1 I142 ( .B(out_70), .A(out_142), .Z(net_142) );
nand2x1 I143 ( .B(out_71), .A(out_143), .Z(net_143) );
nand2x1 I144 ( .B(out_71), .A(out_144), .Z(net_144) );
nand2x1 I145 ( .B(out_72), .A(out_145), .Z(net_145) );
nand2x1 I146 ( .B(out_72), .A(out_146), .Z(net_146) );
nand2x1 I147 ( .B(out_73), .A(out_147), .Z(net_147) );
nand2x1 I148 ( .B(out_73), .A(out_148), .Z(net_148) );
nand2x1 I149 ( .B(out_74), .A(out_149), .Z(net_149) );
nand2x1 I150 ( .B(out_74), .A(out_150), .Z(net_150) );
nand2x1 I151 ( .B(out_75), .A(out_151), .Z(net_151) );
nand2x1 I152 ( .B(out_75), .A(out_152), .Z(net_152) );
nand2x1 I153 ( .B(out_76), .A(out_153), .Z(net_153) );
nand2x1 I154 ( .B(out_76), .A(out_154), .Z(net_154) );
nand2x1 I155 ( .B(out_77), .A(out_155), .Z(net_155) );
nand2x1 I156 ( .B(out_77), .A(out_156), .Z(net_156) );
nand2x1 I157 ( .B(out_78), .A(out_157), .Z(net_157) );
nand2x1 I158 ( .B(out_78), .A(out_158), .Z(net_158) );
nand2x1 I159 ( .B(out_79), .A(out_159), .Z(net_159) );
nand2x1 I160 ( .B(out_79), .A(out_160), .Z(net_160) );
nand2x1 I161 ( .B(out_80), .A(out_161), .Z(net_161) );
nand2x1 I162 ( .B(out_80), .A(out_162), .Z(net_162) );
nand2x1 I163 ( .B(out_81), .A(out_163), .Z(net_163) );
nand2x1 I164 ( .B(out_81), .A(out_164), .Z(net_164) );
nand2x1 I165 ( .B(out_82), .A(out_165), .Z(net_165) );
nand2x1 I166 ( .B(out_82), .A(out_166), .Z(net_166) );
nand2x1 I167 ( .B(out_83), .A(out_167), .Z(net_167) );
nand2x1 I168 ( .B(out_83), .A(out_168), .Z(net_168) );
nand2x1 I169 ( .B(out_84), .A(out_169), .Z(net_169) );
nand2x1 I170 ( .B(out_84), .A(out_170), .Z(net_170) );
nand2x1 I171 ( .B(out_85), .A(out_171), .Z(net_171) );
nand2x1 I172 ( .B(out_85), .A(out_172), .Z(net_172) );
nand2x1 I173 ( .B(out_86), .A(out_173), .Z(net_173) );
nand2x1 I174 ( .B(out_86), .A(out_174), .Z(net_174) );
nand2x1 I175 ( .B(out_87), .A(out_175), .Z(net_175) );
nand2x1 I176 ( .B(out_87), .A(out_176), .Z(net_176) );
nand2x1 I177 ( .B(out_88), .A(out_177), .Z(net_177) );
nand2x1 I178 ( .B(out_88), .A(out_178), .Z(net_178) );
nand2x1 I179 ( .B(out_89), .A(out_179), .Z(net_179) );
nand2x1 I180 ( .B(out_89), .A(out_180), .Z(net_180) );
nand2x1 I181 ( .B(out_90), .A(out_181), .Z(net_181) );
nand2x1 I182 ( .B(out_90), .A(out_182), .Z(net_182) );
nand2x1 I183 ( .B(out_91), .A(out_183), .Z(net_183) );
nand2x1 I184 ( .B(out_91), .A(out_184), .Z(net_184) );
nand2x1 I185 ( .B(out_92), .A(out_185), .Z(net_185) );
nand2x1 I186 ( .B(out_92), .A(out_186), .Z(net_186) );
nand2x1 I187 ( .B(out_93), .A(out_187), .Z(net_187) );
nand2x1 I188 ( .B(out_93), .A(out_188), .Z(net_188) );
nand2x1 I189 ( .B(out_94), .A(out_189), .Z(net_189) );
nand2x1 I190 ( .B(out_94), .A(out_190), .Z(net_190) );
nand2x1 I191 ( .B(out_95), .A(out_191), .Z(net_191) );
nand2x1 I192 ( .B(out_95), .A(out_192), .Z(net_192) );
nand2x1 I193 ( .B(out_96), .A(out_193), .Z(net_193) );
nand2x1 I194 ( .B(out_96), .A(out_194), .Z(net_194) );
nand2x1 I195 ( .B(out_97), .A(out_195), .Z(net_195) );
nand2x1 I196 ( .B(out_97), .A(out_196), .Z(net_196) );
nand2x1 I197 ( .B(out_98), .A(out_197), .Z(net_197) );
nand2x1 I198 ( .B(out_98), .A(out_198), .Z(net_198) );
nand2x1 I199 ( .B(out_99), .A(out_199), .Z(net_199) );
nand2x1 I200 ( .B(out_99), .A(out_200), .Z(net_200) );
nand2x1 I201 ( .B(out_100), .A(out_201), .Z(net_201) );
nand2x1 I202 ( .B(out_100), .A(out_202), .Z(net_202) );
nand2x1 I203 ( .B(out_101), .A(out_203), .Z(net_203) );
nand2x1 I204 ( .B(out_101), .A(out_204), .Z(net_204) );
nand2x1 I205 ( .B(out_102), .A(out_205), .Z(net_205) );
nand2x1 I206 ( .B(out_102), .A(out_206), .Z(net_206) );
nand2x1 I207 ( .B(out_103), .A(out_207), .Z(net_207) );
nand2x1 I208 ( .B(out_103), .A(out_208), .Z(net_208) );
nand2x1 I209 ( .B(out_104), .A(out_209), .Z(net_209) );
nand2x1 I210 ( .B(out_104), .A(out_210), .Z(net_210) );
nand2x1 I211 ( .B(out_105), .A(out_211), .Z(net_211) );
nand2x1 I212 ( .B(out_105), .A(out_212), .Z(net_212) );
nand2x1 I213 ( .B(out_106), .A(out_213), .Z(net_213) );
nand2x1 I214 ( .B(out_106), .A(out_214), .Z(net_214) );
nand2x1 I215 ( .B(out_107), .A(out_215), .Z(net_215) );
nand2x1 I216 ( .B(out_107), .A(out_216), .Z(net_216) );
nand2x1 I217 ( .B(out_108), .A(out_217), .Z(net_217) );
nand2x1 I218 ( .B(out_108), .A(out_218), .Z(net_218) );
nand2x1 I219 ( .B(out_109), .A(out_219), .Z(net_219) );
nand2x1 I220 ( .B(out_109), .A(out_220), .Z(net_220) );
nand2x1 I221 ( .B(out_110), .A(out_221), .Z(net_221) );
nand2x1 I222 ( .B(out_110), .A(out_222), .Z(net_222) );
nand2x1 I223 ( .B(out_111), .A(out_223), .Z(net_223) );
nand2x1 I224 ( .B(out_111), .A(out_224), .Z(net_224) );
nand2x1 I225 ( .B(out_112), .A(out_225), .Z(net_225) );
nand2x1 I226 ( .B(out_112), .A(out_226), .Z(net_226) );
nand2x1 I227 ( .B(out_113), .A(out_227), .Z(net_227) );
nand2x1 I228 ( .B(out_113), .A(out_228), .Z(net_228) );
nand2x1 I229 ( .B(out_114), .A(out_229), .Z(net_229) );
nand2x1 I230 ( .B(out_114), .A(out_230), .Z(net_230) );
nand2x1 I231 ( .B(out_115), .A(out_231), .Z(net_231) );
nand2x1 I232 ( .B(out_115), .A(out_232), .Z(net_232) );
nand2x1 I233 ( .B(out_116), .A(out_233), .Z(net_233) );
nand2x1 I234 ( .B(out_116), .A(out_234), .Z(net_234) );
nand2x1 I235 ( .B(out_117), .A(out_235), .Z(net_235) );
nand2x1 I236 ( .B(out_117), .A(out_236), .Z(net_236) );
nand2x1 I237 ( .B(out_118), .A(out_237), .Z(net_237) );
nand2x1 I238 ( .B(out_118), .A(out_238), .Z(net_238) );
nand2x1 I239 ( .B(out_119), .A(out_239), .Z(net_239) );
nand2x1 I240 ( .B(out_119), .A(out_240), .Z(net_240) );
nand2x1 I241 ( .B(out_120), .A(out_241), .Z(net_241) );
nand2x1 I242 ( .B(out_120), .A(out_242), .Z(net_242) );
nand2x1 I243 ( .B(out_121), .A(out_243), .Z(net_243) );
nand2x1 I244 ( .B(out_121), .A(out_244), .Z(net_244) );
nand2x1 I245 ( .B(out_122), .A(out_245), .Z(net_245) );
nand2x1 I246 ( .B(out_122), .A(out_246), .Z(net_246) );
nand2x1 I247 ( .B(out_123), .A(out_247), .Z(net_247) );
nand2x1 I248 ( .B(out_123), .A(out_248), .Z(net_248) );
nand2x1 I249 ( .B(out_124), .A(out_249), .Z(net_249) );
nand2x1 I250 ( .B(out_124), .A(out_250), .Z(net_250) );
nand2x1 I251 ( .B(out_125), .A(out_251), .Z(net_251) );
nand2x1 I252 ( .B(out_125), .A(out_252), .Z(net_252) );
nand2x1 I253 ( .B(out_126), .A(out_253), .Z(net_253) );
nand2x1 I254 ( .B(out_126), .A(out_254), .Z(net_254) );
nand2x1 I255 ( .B(out_127), .A(out_255), .Z(net_255) );
nand2x1 I256 ( .B(out_127), .A(out_256), .Z(net_256) );
nand2x1 I257 ( .B(out_128), .A(out_257), .Z(net_257) );
nand2x1 I258 ( .B(out_128), .A(out_258), .Z(net_258) );
nand2x1 I259 ( .B(out_129), .A(out_259), .Z(net_259) );
nand2x1 I260 ( .B(out_129), .A(out_260), .Z(net_260) );
nand2x1 I261 ( .B(out_130), .A(out_261), .Z(net_261) );
nand2x1 I262 ( .B(out_130), .A(out_262), .Z(net_262) );
nand2x1 I263 ( .B(out_131), .A(out_263), .Z(net_263) );
nand2x1 I264 ( .B(out_131), .A(out_264), .Z(net_264) );
nand2x1 I265 ( .B(out_132), .A(out_265), .Z(net_265) );
nand2x1 I266 ( .B(out_132), .A(out_266), .Z(net_266) );
endmodule
